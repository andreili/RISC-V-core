@0
00000033
40000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
