@0
00000033
00100093
40000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
00000033
